
`timescale 1ns / 1ps


//Clk??????????
//Reset??????????
//Result????????????????????????????
//Addr??????????
module PC(Clk,Reset,Result,Address);  
input Clk;//??
input Reset;//????PC??????     
input[31:0] Result;
output reg[31:0] Address;

//address ????0
initial begin
Address  <= 0;
end

always @(posedge Clk or negedge Reset)  //
begin  
if (!Reset) //????????????address??0
	begin  
	Address <= 0;  
	end  
else   
	begin
	Address =  Result; //????pc? 
	end  
end  
endmodule


//??32???????pc?4???
module PCadd4(PC_o,PCadd4);
input [31:0] PC_o;//???
output [31:0] PCadd4;//?????
CLA_32 cla32(PC_o,4,0, PCadd4, Cout);

endmodule
