module ORgate(in1,in2,Out);

input in1,in2;
output Out;

assign Out=in1|in2;

endmodule

